
package barrel_shifter_pkg;
    parameter int WIDTH = 8;
endpackage
