
package fifo_buffer_pkg;
    parameter int DATA_WIDTH    = 8;
    parameter int DEPTH         = 16;
endpackage
