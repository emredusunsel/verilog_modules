
package clock_divider_pkg;
    parameter int DIV = 2;
endpackage
