
package fwft_fifo_pkg;
    parameter int DATA_WIDTH    = 32;
    parameter int DEPTH         = 16;
endpackage
