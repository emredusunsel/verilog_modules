
package onehot_to_binary_pkg;
    parameter int STATE_W   = 8;
    parameter int BIN_W     = $clog2(STATE_W);
endpackage
