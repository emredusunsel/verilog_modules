
package mux_pkg;
    parameter int   WIDTH   = 32;
    parameter int   N       = 4;
endpackage
