
package register_file_pkg;
    parameter int DATA_WIDTH    = 32;
    parameter int REG_COUNT     = 8;
    parameter int ADDR_WIDTH    = $clog2(REG_COUNT);
endpackage
