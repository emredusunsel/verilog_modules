
package register_file_pkg;
    parameter int DATA_WIDTH    = 32;
    parameter int ADDR_WIDTH    = 4;
    parameter int REG_COUNT     = 8;
endpackage
