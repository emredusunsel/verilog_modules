
package counter_pkg;
    parameter int WIDTH = 4;
    typedef enum logic {DOWN=1'b0, UP=1'b1} count_dir_e;
endpackage
