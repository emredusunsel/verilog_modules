
package comparator_pkg;
    parameter int WIDTH = 8;
endpackage
